* C:\Users\naiar\OneDrive\Documentos\NAIARA\ESTUDIO\TCO\pract\pract7\pract7.2.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 16 21:05:06 2020



** Analysis setup **
.tran 0ns 1u
.OP 
.LIB "C:\Users\naiar\OneDrive\Documentos\NAIARA\ESTUDIO\TCO\pract\pract7\pract7.1.lib"
.STMLIB "pract7.2.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "pract7.2.net"
.INC "pract7.2.als"


.probe


.END
