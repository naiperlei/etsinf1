* C:\Users\naiar\OneDrive\Documentos\NAIARA\ESTUDIO\TCO\pract\pract5\pract5.2.sch

* Schematics Version 9.1 - Web Update 1
* Sat May 16 17:32:25 2020



** Analysis setup **
.tran 1n 120n
.OP 
.LIB "C:\Users\naiar\OneDrive\Documentos\NAIARA\ESTUDIO\TCO\pract\pract4\pract4.1.lib"
.LIB "C:\Users\naiar\OneDrive\Documentos\NAIARA\ESTUDIO\TCO\pract\pract5\pract5.1.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "pract5.2.net"
.INC "pract5.2.als"


.probe


.END
